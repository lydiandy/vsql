module test

pub fn test_inert() {
}

pub fn test_update() {
}

pub fn test_delete() {
}
