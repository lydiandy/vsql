module vsql

pub fn (db DB) up() {
	
}

pub fn(db DB) down() {
	
}