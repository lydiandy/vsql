module vsql

pub fn logger() {
	
}