module test

pub fn test_inert() {
	db := connect_db()
	// start to test
	mut res := ''
}

pub fn test_update() {
	db := connect_db()
	// start to test
	mut res := ''
}

pub fn test_delete() {
	db := connect_db()
	// start to test
	mut res := ''
}
