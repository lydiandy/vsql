module test

fn test_schema() {
	db := connect_db()
	// start to test
	mut res := ''
}
