module vsql

pub fn (mut db DB) up() {
}

pub fn (mut db DB) down() {
}
