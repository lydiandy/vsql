module test

fn test_transaction() {
	db := connect_db()
	// start to test
	mut res := ''
}
